package Test;
import Prelude::*;

(* synthesize *)
module mkTest (Empty);
endmodule
endpackage
